library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use std.textio.all;

entity instructionMemory is
    Port ( 
			  --clk : in STD_LOGIC;
			  address : in  STD_LOGIC_VECTOR (31 downto 0);
           reset : in  STD_LOGIC;
           outInstruction : out  STD_LOGIC_VECTOR (31 downto 0));
end instructionMemory;
architecture Behavioral of instructionMemory is

type rom_type is array (63 downto 0) of std_logic_vector (31 downto 0);
signal ROM : rom_type := (	"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
																					-- 6
									"01111111111111111111111111110001", "10100110000100000010000000000110",
									-- 5
									"10100100000100000010000000000101", "00000001000000000000000000000000",
									
									"10000011110000111110000000000000", "10010000000100000000000000010000",
									"00000110101111111111111111111011", "10000000101001000100000000010011",
									"10100010000100000000000000010100", "10101000000001000110000000000001",
									"10100000000100000000000000010100", "10101000000001000000000000010010",
									"00110110100000000000000000001000", "10000000101001000100000000010011",	
									"10100010000100000010000000000000", "10100000000100000010000000000000");

begin

    process (reset,address,ROM)
    begin
        if (reset='1') then
				outInstruction <= "00000000000000000000000000000000";
		  else
            outInstruction <= ROM(conv_integer(address(5 downto 0)));  
        end if;
    end process;
end Behavioral;

